/*
Author: Ian Gilman
Title: 32-bit Set Less Than
Summary: Sets result to 1 if if operand0 is less than operand1 for signed value
   else sets to 0.
*/

module slt(operand0, operand1, result)
   input [31:0] operand0, operand1;
   output [31:0] result;
   
   /* use subtract to solve */
   

endmodule