/*
Author: Ian Gilman
Title: Negate a signed number
Summary: Return the negative value of a signed number
*/

module negate_signed_gate(orig_num, neg_num);
// I/O
   input wire [31:0] orig_num;
   output wire [31:0] neg_num;
// Internal
   
   
   
endmodule